-- calculates roundkeys from cipher (conducts xor operations) 


-- output: 11 128-bit arrays