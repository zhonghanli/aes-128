LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;
USE WORK.aes_const.all;


entity key_init is


end entity key_init;


architecture behavior of key_init is
	TYPE state is (s0,s1,s2);
	signal 

begin

end architecture behavior;